VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_logo
  CLASS BLOCK ;
  FOREIGN skullfet_logo ;
  ORIGIN -50.000 -50.000 ;
  SIZE 700.000 BY 800.000 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 725.000 50.000 750.000 850.000 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 50.000 50.000 75.000 850.000 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 351.500 807.500 459.500 821.000 ;
        RECT 338.000 794.000 459.500 807.500 ;
        RECT 311.000 767.000 486.500 794.000 ;
        RECT 297.500 713.000 500.000 767.000 ;
        RECT 297.500 699.500 338.000 713.000 ;
        RECT 297.500 686.000 324.500 699.500 ;
        RECT 311.000 672.500 324.500 686.000 ;
        RECT 378.500 672.500 419.000 713.000 ;
        RECT 459.500 699.500 500.000 713.000 ;
        RECT 473.000 686.000 500.000 699.500 ;
        RECT 473.000 672.500 486.500 686.000 ;
        RECT 311.000 659.000 338.000 672.500 ;
        RECT 365.000 659.000 432.500 672.500 ;
        RECT 459.500 659.000 486.500 672.500 ;
        RECT 311.000 645.500 392.000 659.000 ;
        RECT 405.500 645.500 473.000 659.000 ;
        RECT 338.000 632.000 378.500 645.500 ;
        RECT 419.000 632.000 473.000 645.500 ;
        RECT 351.500 605.000 446.000 632.000 ;
        RECT 270.500 591.500 311.000 605.000 ;
        RECT 351.500 591.500 365.000 605.000 ;
        RECT 378.500 591.500 392.000 605.000 ;
        RECT 405.500 591.500 419.000 605.000 ;
        RECT 432.500 591.500 446.000 605.000 ;
        RECT 486.500 591.500 527.000 605.000 ;
        RECT 257.000 564.500 324.500 591.500 ;
        RECT 473.000 564.500 540.500 591.500 ;
        RECT 270.500 551.000 351.500 564.500 ;
        RECT 446.000 551.000 527.000 564.500 ;
        RECT 311.000 537.500 365.000 551.000 ;
        RECT 432.500 537.500 486.500 551.000 ;
        RECT 338.000 524.000 392.000 537.500 ;
        RECT 405.500 524.000 459.500 537.500 ;
        RECT 365.000 497.000 432.500 524.000 ;
        RECT 338.000 483.500 392.000 497.000 ;
        RECT 405.500 483.500 459.500 497.000 ;
        RECT 270.500 470.000 365.000 483.500 ;
        RECT 432.500 470.000 540.500 483.500 ;
        RECT 257.000 456.500 338.000 470.000 ;
        RECT 459.500 456.500 540.500 470.000 ;
        RECT 257.000 443.000 311.000 456.500 ;
        RECT 486.500 443.000 540.500 456.500 ;
        RECT 257.000 429.500 297.500 443.000 ;
        RECT 500.000 429.500 540.500 443.000 ;
        RECT 270.500 416.000 284.000 429.500 ;
        RECT 351.500 416.000 365.000 429.500 ;
        RECT 378.500 416.000 392.000 429.500 ;
        RECT 405.500 416.000 419.000 429.500 ;
        RECT 432.500 416.000 446.000 429.500 ;
        RECT 513.500 416.000 527.000 429.500 ;
        RECT 351.500 389.000 446.000 416.000 ;
        RECT 338.000 375.500 378.500 389.000 ;
        RECT 419.000 375.500 473.000 389.000 ;
        RECT 311.000 362.000 392.000 375.500 ;
        RECT 405.500 362.000 473.000 375.500 ;
        RECT 311.000 348.500 338.000 362.000 ;
        RECT 365.000 348.500 432.500 362.000 ;
        RECT 459.500 348.500 486.500 362.000 ;
        RECT 311.000 335.000 324.500 348.500 ;
        RECT 297.500 321.500 324.500 335.000 ;
        RECT 297.500 308.000 338.000 321.500 ;
        RECT 378.500 308.000 419.000 348.500 ;
        RECT 473.000 335.000 486.500 348.500 ;
        RECT 473.000 321.500 500.000 335.000 ;
        RECT 459.500 308.000 500.000 321.500 ;
        RECT 297.500 254.000 500.000 308.000 ;
        RECT 311.000 227.000 486.500 254.000 ;
        RECT 338.000 213.500 459.500 227.000 ;
        RECT 351.500 200.000 459.500 213.500 ;
        RECT 170.000 155.000 210.000 160.000 ;
        RECT 235.000 155.000 240.000 160.000 ;
        RECT 260.000 155.000 265.000 160.000 ;
        RECT 165.000 150.000 210.000 155.000 ;
        RECT 230.000 150.000 240.000 155.000 ;
        RECT 255.000 150.000 270.000 155.000 ;
        RECT 160.000 120.000 175.000 150.000 ;
        RECT 195.000 140.000 210.000 150.000 ;
        RECT 195.000 135.000 205.000 140.000 ;
        RECT 195.000 130.000 200.000 135.000 ;
        RECT 225.000 130.000 240.000 150.000 ;
        RECT 250.000 145.000 270.000 150.000 ;
        RECT 245.000 140.000 265.000 145.000 ;
        RECT 245.000 135.000 260.000 140.000 ;
        RECT 245.000 130.000 255.000 135.000 ;
        RECT 225.000 125.000 255.000 130.000 ;
        RECT 220.000 120.000 250.000 125.000 ;
        RECT 150.000 115.000 210.000 120.000 ;
        RECT 215.000 115.000 250.000 120.000 ;
        RECT 155.000 110.000 210.000 115.000 ;
        RECT 170.000 95.000 175.000 100.000 ;
        RECT 165.000 90.000 175.000 95.000 ;
        RECT 195.000 90.000 210.000 110.000 ;
        RECT 225.000 110.000 255.000 115.000 ;
        RECT 160.000 85.000 205.000 90.000 ;
        RECT 155.000 80.000 200.000 85.000 ;
        RECT 225.000 80.000 240.000 110.000 ;
        RECT 245.000 105.000 255.000 110.000 ;
        RECT 245.000 100.000 260.000 105.000 ;
        RECT 245.000 95.000 265.000 100.000 ;
        RECT 250.000 90.000 270.000 95.000 ;
        RECT 255.000 85.000 270.000 90.000 ;
        RECT 275.000 90.000 290.000 160.000 ;
        RECT 310.000 155.000 315.000 160.000 ;
        RECT 340.000 155.000 345.000 160.000 ;
        RECT 390.000 155.000 395.000 160.000 ;
        RECT 450.000 155.000 490.000 160.000 ;
        RECT 515.000 155.000 555.000 160.000 ;
        RECT 310.000 150.000 320.000 155.000 ;
        RECT 335.000 150.000 345.000 155.000 ;
        RECT 385.000 150.000 395.000 155.000 ;
        RECT 445.000 150.000 490.000 155.000 ;
        RECT 510.000 150.000 555.000 155.000 ;
        RECT 580.000 150.000 595.000 160.000 ;
        RECT 310.000 90.000 325.000 150.000 ;
        RECT 330.000 90.000 345.000 150.000 ;
        RECT 370.000 90.000 375.000 95.000 ;
        RECT 275.000 85.000 320.000 90.000 ;
        RECT 330.000 85.000 355.000 90.000 ;
        RECT 365.000 85.000 375.000 90.000 ;
        RECT 260.000 80.000 265.000 85.000 ;
        RECT 275.000 80.000 315.000 85.000 ;
        RECT 330.000 80.000 375.000 85.000 ;
        RECT 380.000 90.000 395.000 150.000 ;
        RECT 440.000 125.000 455.000 150.000 ;
        RECT 475.000 140.000 490.000 150.000 ;
        RECT 475.000 135.000 485.000 140.000 ;
        RECT 475.000 130.000 480.000 135.000 ;
        RECT 505.000 125.000 520.000 150.000 ;
        RECT 540.000 140.000 555.000 150.000 ;
        RECT 560.000 145.000 610.000 150.000 ;
        RECT 565.000 140.000 615.000 145.000 ;
        RECT 540.000 135.000 550.000 140.000 ;
        RECT 575.000 135.000 615.000 140.000 ;
        RECT 540.000 130.000 545.000 135.000 ;
        RECT 435.000 120.000 470.000 125.000 ;
        RECT 500.000 120.000 535.000 125.000 ;
        RECT 430.000 115.000 470.000 120.000 ;
        RECT 495.000 115.000 535.000 120.000 ;
        RECT 420.000 90.000 425.000 95.000 ;
        RECT 380.000 85.000 405.000 90.000 ;
        RECT 415.000 85.000 425.000 90.000 ;
        RECT 380.000 80.000 425.000 85.000 ;
        RECT 440.000 80.000 455.000 115.000 ;
        RECT 505.000 90.000 520.000 115.000 ;
        RECT 540.000 105.000 545.000 110.000 ;
        RECT 540.000 100.000 550.000 105.000 ;
        RECT 540.000 90.000 555.000 100.000 ;
        RECT 505.000 80.000 555.000 90.000 ;
        RECT 580.000 90.000 595.000 135.000 ;
        RECT 605.000 130.000 615.000 135.000 ;
        RECT 610.000 125.000 615.000 130.000 ;
        RECT 580.000 85.000 605.000 90.000 ;
        RECT 575.000 80.000 600.000 85.000 ;
        RECT 225.000 75.000 230.000 80.000 ;
        RECT 330.000 75.000 335.000 80.000 ;
        RECT 380.000 75.000 385.000 80.000 ;
      LAYER Metal2 ;
        RECT 250.000 200.000 550.000 850.000 ;
        RECT 125.000 50.000 650.000 200.000 ;
      LAYER Metal3 ;
        RECT 250.000 200.000 550.000 850.000 ;
        RECT 125.000 50.000 650.000 200.000 ;
      LAYER Metal4 ;
        RECT 351.500 807.500 459.500 821.000 ;
        RECT 338.000 794.000 459.500 807.500 ;
        RECT 311.000 767.000 486.500 794.000 ;
        RECT 297.500 713.000 500.000 767.000 ;
        RECT 297.500 699.500 338.000 713.000 ;
        RECT 297.500 686.000 324.500 699.500 ;
        RECT 311.000 672.500 324.500 686.000 ;
        RECT 378.500 672.500 419.000 713.000 ;
        RECT 459.500 699.500 500.000 713.000 ;
        RECT 473.000 686.000 500.000 699.500 ;
        RECT 473.000 672.500 486.500 686.000 ;
        RECT 311.000 659.000 338.000 672.500 ;
        RECT 365.000 659.000 432.500 672.500 ;
        RECT 459.500 659.000 486.500 672.500 ;
        RECT 311.000 645.500 392.000 659.000 ;
        RECT 405.500 645.500 473.000 659.000 ;
        RECT 338.000 632.000 378.500 645.500 ;
        RECT 419.000 632.000 473.000 645.500 ;
        RECT 351.500 605.000 446.000 632.000 ;
        RECT 270.500 591.500 311.000 605.000 ;
        RECT 351.500 591.500 365.000 605.000 ;
        RECT 378.500 591.500 392.000 605.000 ;
        RECT 405.500 591.500 419.000 605.000 ;
        RECT 432.500 591.500 446.000 605.000 ;
        RECT 486.500 591.500 527.000 605.000 ;
        RECT 257.000 564.500 324.500 591.500 ;
        RECT 473.000 564.500 540.500 591.500 ;
        RECT 270.500 551.000 351.500 564.500 ;
        RECT 446.000 551.000 527.000 564.500 ;
        RECT 311.000 537.500 365.000 551.000 ;
        RECT 432.500 537.500 486.500 551.000 ;
        RECT 338.000 524.000 392.000 537.500 ;
        RECT 405.500 524.000 459.500 537.500 ;
        RECT 365.000 497.000 432.500 524.000 ;
        RECT 338.000 483.500 392.000 497.000 ;
        RECT 405.500 483.500 459.500 497.000 ;
        RECT 270.500 470.000 365.000 483.500 ;
        RECT 432.500 470.000 540.500 483.500 ;
        RECT 257.000 456.500 338.000 470.000 ;
        RECT 459.500 456.500 540.500 470.000 ;
        RECT 257.000 443.000 311.000 456.500 ;
        RECT 486.500 443.000 540.500 456.500 ;
        RECT 257.000 429.500 297.500 443.000 ;
        RECT 500.000 429.500 540.500 443.000 ;
        RECT 270.500 416.000 284.000 429.500 ;
        RECT 351.500 416.000 365.000 429.500 ;
        RECT 378.500 416.000 392.000 429.500 ;
        RECT 405.500 416.000 419.000 429.500 ;
        RECT 432.500 416.000 446.000 429.500 ;
        RECT 513.500 416.000 527.000 429.500 ;
        RECT 351.500 389.000 446.000 416.000 ;
        RECT 338.000 375.500 378.500 389.000 ;
        RECT 419.000 375.500 473.000 389.000 ;
        RECT 311.000 362.000 392.000 375.500 ;
        RECT 405.500 362.000 473.000 375.500 ;
        RECT 311.000 348.500 338.000 362.000 ;
        RECT 365.000 348.500 432.500 362.000 ;
        RECT 459.500 348.500 486.500 362.000 ;
        RECT 311.000 335.000 324.500 348.500 ;
        RECT 297.500 321.500 324.500 335.000 ;
        RECT 297.500 308.000 338.000 321.500 ;
        RECT 378.500 308.000 419.000 348.500 ;
        RECT 473.000 335.000 486.500 348.500 ;
        RECT 473.000 321.500 500.000 335.000 ;
        RECT 459.500 308.000 500.000 321.500 ;
        RECT 297.500 254.000 500.000 308.000 ;
        RECT 311.000 227.000 486.500 254.000 ;
        RECT 338.000 213.500 459.500 227.000 ;
        RECT 351.500 200.000 459.500 213.500 ;
        RECT 170.000 155.000 210.000 160.000 ;
        RECT 235.000 155.000 240.000 160.000 ;
        RECT 260.000 155.000 265.000 160.000 ;
        RECT 165.000 150.000 210.000 155.000 ;
        RECT 230.000 150.000 240.000 155.000 ;
        RECT 255.000 150.000 270.000 155.000 ;
        RECT 160.000 120.000 175.000 150.000 ;
        RECT 195.000 140.000 210.000 150.000 ;
        RECT 195.000 135.000 205.000 140.000 ;
        RECT 195.000 130.000 200.000 135.000 ;
        RECT 225.000 130.000 240.000 150.000 ;
        RECT 250.000 145.000 270.000 150.000 ;
        RECT 245.000 140.000 265.000 145.000 ;
        RECT 245.000 135.000 260.000 140.000 ;
        RECT 245.000 130.000 255.000 135.000 ;
        RECT 225.000 125.000 255.000 130.000 ;
        RECT 220.000 120.000 250.000 125.000 ;
        RECT 150.000 115.000 210.000 120.000 ;
        RECT 215.000 115.000 250.000 120.000 ;
        RECT 155.000 110.000 210.000 115.000 ;
        RECT 170.000 95.000 175.000 100.000 ;
        RECT 165.000 90.000 175.000 95.000 ;
        RECT 195.000 90.000 210.000 110.000 ;
        RECT 225.000 110.000 255.000 115.000 ;
        RECT 160.000 85.000 205.000 90.000 ;
        RECT 155.000 80.000 200.000 85.000 ;
        RECT 225.000 80.000 240.000 110.000 ;
        RECT 245.000 105.000 255.000 110.000 ;
        RECT 245.000 100.000 260.000 105.000 ;
        RECT 245.000 95.000 265.000 100.000 ;
        RECT 250.000 90.000 270.000 95.000 ;
        RECT 255.000 85.000 270.000 90.000 ;
        RECT 275.000 90.000 290.000 160.000 ;
        RECT 310.000 155.000 315.000 160.000 ;
        RECT 340.000 155.000 345.000 160.000 ;
        RECT 390.000 155.000 395.000 160.000 ;
        RECT 450.000 155.000 490.000 160.000 ;
        RECT 515.000 155.000 555.000 160.000 ;
        RECT 310.000 150.000 320.000 155.000 ;
        RECT 335.000 150.000 345.000 155.000 ;
        RECT 385.000 150.000 395.000 155.000 ;
        RECT 445.000 150.000 490.000 155.000 ;
        RECT 510.000 150.000 555.000 155.000 ;
        RECT 580.000 150.000 595.000 160.000 ;
        RECT 310.000 90.000 325.000 150.000 ;
        RECT 330.000 90.000 345.000 150.000 ;
        RECT 370.000 90.000 375.000 95.000 ;
        RECT 275.000 85.000 320.000 90.000 ;
        RECT 330.000 85.000 355.000 90.000 ;
        RECT 365.000 85.000 375.000 90.000 ;
        RECT 260.000 80.000 265.000 85.000 ;
        RECT 275.000 80.000 315.000 85.000 ;
        RECT 330.000 80.000 375.000 85.000 ;
        RECT 380.000 90.000 395.000 150.000 ;
        RECT 440.000 125.000 455.000 150.000 ;
        RECT 475.000 140.000 490.000 150.000 ;
        RECT 475.000 135.000 485.000 140.000 ;
        RECT 475.000 130.000 480.000 135.000 ;
        RECT 505.000 125.000 520.000 150.000 ;
        RECT 540.000 140.000 555.000 150.000 ;
        RECT 560.000 145.000 610.000 150.000 ;
        RECT 565.000 140.000 615.000 145.000 ;
        RECT 540.000 135.000 550.000 140.000 ;
        RECT 575.000 135.000 615.000 140.000 ;
        RECT 540.000 130.000 545.000 135.000 ;
        RECT 435.000 120.000 470.000 125.000 ;
        RECT 500.000 120.000 535.000 125.000 ;
        RECT 430.000 115.000 470.000 120.000 ;
        RECT 495.000 115.000 535.000 120.000 ;
        RECT 420.000 90.000 425.000 95.000 ;
        RECT 380.000 85.000 405.000 90.000 ;
        RECT 415.000 85.000 425.000 90.000 ;
        RECT 380.000 80.000 425.000 85.000 ;
        RECT 440.000 80.000 455.000 115.000 ;
        RECT 505.000 90.000 520.000 115.000 ;
        RECT 540.000 105.000 545.000 110.000 ;
        RECT 540.000 100.000 550.000 105.000 ;
        RECT 540.000 90.000 555.000 100.000 ;
        RECT 505.000 80.000 555.000 90.000 ;
        RECT 580.000 90.000 595.000 135.000 ;
        RECT 605.000 130.000 615.000 135.000 ;
        RECT 610.000 125.000 615.000 130.000 ;
        RECT 580.000 85.000 605.000 90.000 ;
        RECT 575.000 80.000 600.000 85.000 ;
        RECT 225.000 75.000 230.000 80.000 ;
        RECT 330.000 75.000 335.000 80.000 ;
        RECT 380.000 75.000 385.000 80.000 ;
  END
END skullfet_logo
END LIBRARY

