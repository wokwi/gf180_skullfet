VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_nand
  CLASS BLOCK ;
  FOREIGN skullfet_nand ;
  ORIGIN 0.000 -5.400 ;
  SIZE 81.000 BY 66.150 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 109.349998 ;
    PORT
      LAYER Metal1 ;
        RECT 58.725 60.075 72.225 62.775 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 109.349998 ;
    PORT
      LAYER Metal1 ;
        RECT 8.775 14.175 22.275 16.875 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 442.867493 ;
    PORT
      LAYER Metal1 ;
        RECT 47.925 56.700 57.375 59.400 ;
        RECT 54.675 54.000 68.850 56.700 ;
        RECT 66.150 46.575 68.850 54.000 ;
        RECT 66.150 20.250 68.850 31.725 ;
        RECT 47.925 17.550 68.850 20.250 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 73.575 12.825 76.275 33.075 ;
        RECT 46.575 10.125 76.275 12.825 ;
      LAYER Via1 ;
        RECT 74.250 10.800 75.600 12.150 ;
      LAYER Metal2 ;
        RECT 73.575 10.125 76.275 12.825 ;
      LAYER Via2 ;
        RECT 74.250 10.800 75.600 12.150 ;
      LAYER Metal3 ;
        RECT 73.575 10.125 76.275 12.825 ;
      LAYER Via3 ;
        RECT 74.250 10.800 75.600 12.150 ;
      LAYER Metal4 ;
        RECT 73.575 5.400 76.275 71.550 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.725 5.400 7.425 33.075 ;
      LAYER Via1 ;
        RECT 5.400 27.675 6.750 29.025 ;
      LAYER Metal2 ;
        RECT 7.425 47.925 15.525 49.275 ;
        RECT 4.725 46.575 18.225 47.925 ;
        RECT 4.725 45.225 14.175 46.575 ;
        RECT 16.875 45.225 20.925 46.575 ;
        RECT 2.025 41.175 12.825 45.225 ;
        RECT 18.225 43.875 20.925 45.225 ;
        RECT 18.225 42.525 24.975 43.875 ;
        RECT 16.875 41.175 23.625 42.525 ;
        RECT 2.025 39.825 19.575 41.175 ;
        RECT 20.925 39.825 24.975 41.175 ;
        RECT 2.025 38.475 18.225 39.825 ;
        RECT 20.925 38.475 23.625 39.825 ;
        RECT 2.025 37.125 19.575 38.475 ;
        RECT 20.925 37.125 24.975 38.475 ;
        RECT 2.025 34.425 12.825 37.125 ;
        RECT 16.875 35.775 23.625 37.125 ;
        RECT 3.375 33.075 12.825 34.425 ;
        RECT 18.225 34.425 24.975 35.775 ;
        RECT 18.225 33.075 20.925 34.425 ;
        RECT 4.725 31.725 14.175 33.075 ;
        RECT 16.875 31.725 19.575 33.075 ;
        RECT 4.725 30.375 19.575 31.725 ;
        RECT 7.425 29.700 15.525 30.375 ;
        RECT 4.725 29.025 15.525 29.700 ;
        RECT 4.725 27.000 7.425 29.025 ;
      LAYER Via2 ;
        RECT 5.400 27.675 6.750 29.025 ;
      LAYER Metal3 ;
        RECT 4.725 27.000 7.425 29.700 ;
      LAYER Via3 ;
        RECT 5.400 27.675 6.750 29.025 ;
      LAYER Metal4 ;
        RECT 4.725 5.400 7.425 71.550 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 12.150 64.125 34.425 66.825 ;
        RECT 12.150 46.575 14.850 64.125 ;
        RECT 27.675 46.575 30.375 47.925 ;
        RECT 50.625 46.575 53.325 47.925 ;
        RECT 26.325 43.875 33.075 46.575 ;
        RECT 47.925 43.875 54.675 46.575 ;
        RECT 27.675 42.525 35.775 43.875 ;
        RECT 45.225 42.525 53.325 43.875 ;
        RECT 31.725 41.175 37.125 42.525 ;
        RECT 43.875 41.175 49.275 42.525 ;
        RECT 34.425 39.825 39.825 41.175 ;
        RECT 41.175 39.825 46.575 41.175 ;
        RECT 37.125 37.125 43.875 39.825 ;
        RECT 34.425 35.775 39.825 37.125 ;
        RECT 41.175 35.775 46.575 37.125 ;
        RECT 27.675 34.425 37.125 35.775 ;
        RECT 43.875 34.425 54.675 35.775 ;
        RECT 26.325 33.075 34.425 34.425 ;
        RECT 46.575 33.075 54.675 34.425 ;
        RECT 26.325 31.725 31.725 33.075 ;
        RECT 49.275 31.725 54.675 33.075 ;
        RECT 26.325 30.375 30.375 31.725 ;
        RECT 50.625 30.375 54.675 31.725 ;
        RECT 27.675 29.025 29.025 30.375 ;
        RECT 51.975 29.025 53.325 30.375 ;
      LAYER Metal2 ;
        RECT 35.775 68.175 46.575 69.525 ;
        RECT 34.425 66.825 46.575 68.175 ;
        RECT 31.725 64.125 49.275 66.825 ;
        RECT 30.375 58.725 50.625 64.125 ;
        RECT 30.375 57.375 34.425 58.725 ;
        RECT 30.375 56.025 33.075 57.375 ;
        RECT 31.725 54.675 33.075 56.025 ;
        RECT 38.475 54.675 42.525 58.725 ;
        RECT 46.575 57.375 50.625 58.725 ;
        RECT 47.925 56.025 50.625 57.375 ;
        RECT 47.925 54.675 49.275 56.025 ;
        RECT 31.725 53.325 34.425 54.675 ;
        RECT 37.125 53.325 43.875 54.675 ;
        RECT 46.575 53.325 49.275 54.675 ;
        RECT 31.725 51.975 39.825 53.325 ;
        RECT 41.175 51.975 47.925 53.325 ;
        RECT 34.425 50.625 38.475 51.975 ;
        RECT 42.525 50.625 47.925 51.975 ;
        RECT 35.775 47.925 45.225 50.625 ;
        RECT 65.475 47.925 73.575 49.275 ;
        RECT 35.775 46.575 37.125 47.925 ;
        RECT 38.475 46.575 39.825 47.925 ;
        RECT 41.175 46.575 42.525 47.925 ;
        RECT 43.875 46.575 45.225 47.925 ;
        RECT 61.425 46.575 76.275 47.925 ;
        RECT 61.425 45.225 64.125 46.575 ;
        RECT 66.825 45.225 76.275 46.575 ;
        RECT 60.075 43.875 62.775 45.225 ;
        RECT 56.025 42.525 62.775 43.875 ;
        RECT 68.175 43.875 77.625 45.225 ;
        RECT 57.375 41.175 64.125 42.525 ;
        RECT 68.175 41.175 78.975 43.875 ;
        RECT 56.025 39.825 60.075 41.175 ;
        RECT 61.425 39.825 78.975 41.175 ;
        RECT 57.375 38.475 60.075 39.825 ;
        RECT 62.775 38.475 78.975 39.825 ;
        RECT 56.025 37.125 60.075 38.475 ;
        RECT 61.425 37.125 78.975 38.475 ;
        RECT 57.375 35.775 64.125 37.125 ;
        RECT 56.025 34.425 62.775 35.775 ;
        RECT 60.075 33.075 62.775 34.425 ;
        RECT 68.175 33.075 78.975 37.125 ;
        RECT 60.075 31.725 64.125 33.075 ;
        RECT 66.825 31.725 76.275 33.075 ;
        RECT 62.775 30.375 76.275 31.725 ;
        RECT 35.775 29.025 37.125 30.375 ;
        RECT 38.475 29.025 39.825 30.375 ;
        RECT 41.175 29.025 42.525 30.375 ;
        RECT 43.875 29.025 45.225 30.375 ;
        RECT 65.475 29.025 73.575 30.375 ;
        RECT 35.775 26.325 45.225 29.025 ;
        RECT 34.425 24.975 38.475 26.325 ;
        RECT 42.525 24.975 47.925 26.325 ;
        RECT 31.725 23.625 39.825 24.975 ;
        RECT 41.175 23.625 47.925 24.975 ;
        RECT 31.725 22.275 34.425 23.625 ;
        RECT 37.125 22.275 43.875 23.625 ;
        RECT 46.575 22.275 49.275 23.625 ;
        RECT 31.725 20.925 33.075 22.275 ;
        RECT 30.375 19.575 33.075 20.925 ;
        RECT 30.375 18.225 34.425 19.575 ;
        RECT 38.475 18.225 42.525 22.275 ;
        RECT 47.925 20.925 49.275 22.275 ;
        RECT 47.925 19.575 50.625 20.925 ;
        RECT 46.575 18.225 50.625 19.575 ;
        RECT 30.375 12.825 50.625 18.225 ;
        RECT 31.725 10.125 49.275 12.825 ;
        RECT 34.425 8.775 46.575 10.125 ;
        RECT 35.775 7.425 46.575 8.775 ;
  END
END skullfet_nand
END LIBRARY

