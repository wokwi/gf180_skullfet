VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 53.500 BY 72.000 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 70.000 53.500 72.000 ;
        RECT 12.500 62.000 14.500 70.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 13.000 2.000 15.200 12.000 ;
        RECT 0.000 0.000 53.500 2.000 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 317.519989 ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 55.750 20.000 58.250 ;
        RECT 12.500 17.750 15.000 55.750 ;
        RECT 12.500 15.250 20.500 17.750 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 81.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 42.500 22.750 45.000 49.750 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 16.500 65.250 20.500 69.000 ;
        RECT 15.500 64.750 21.500 65.250 ;
        RECT 15.500 63.500 16.000 64.750 ;
        RECT 17.250 63.500 21.500 64.750 ;
        RECT 15.500 62.750 21.500 63.500 ;
        RECT 17.000 9.750 21.500 10.750 ;
        RECT 17.000 8.750 17.250 9.750 ;
        RECT 18.500 8.750 21.500 9.750 ;
        RECT 17.000 8.250 21.500 8.750 ;
        RECT 16.750 4.750 20.250 8.250 ;
      LAYER Metal2 ;
        RECT 23.650 66.500 34.450 67.850 ;
        RECT 22.300 65.150 34.450 66.500 ;
        RECT 19.600 62.450 37.150 65.150 ;
        RECT 18.250 57.050 38.500 62.450 ;
        RECT 18.250 55.700 22.300 57.050 ;
        RECT 18.250 54.350 20.950 55.700 ;
        RECT 19.600 53.000 20.950 54.350 ;
        RECT 26.350 53.000 30.400 57.050 ;
        RECT 34.450 55.700 38.500 57.050 ;
        RECT 35.800 54.350 38.500 55.700 ;
        RECT 35.800 53.000 37.150 54.350 ;
        RECT 19.600 51.650 22.300 53.000 ;
        RECT 25.000 51.650 31.750 53.000 ;
        RECT 34.450 51.650 37.150 53.000 ;
        RECT 19.600 50.300 27.700 51.650 ;
        RECT 29.050 50.300 35.800 51.650 ;
        RECT 22.300 48.950 26.350 50.300 ;
        RECT 30.400 48.950 35.800 50.300 ;
        RECT 23.650 46.250 33.100 48.950 ;
        RECT 15.550 44.900 19.600 46.250 ;
        RECT 23.650 44.900 25.000 46.250 ;
        RECT 26.350 44.900 27.700 46.250 ;
        RECT 29.050 44.900 30.400 46.250 ;
        RECT 31.750 44.900 33.100 46.250 ;
        RECT 37.150 44.900 41.200 46.250 ;
        RECT 14.200 42.200 20.950 44.900 ;
        RECT 35.800 42.200 42.550 44.900 ;
        RECT 15.550 40.850 23.650 42.200 ;
        RECT 33.100 40.850 41.200 42.200 ;
        RECT 19.600 39.500 25.000 40.850 ;
        RECT 31.750 39.500 37.150 40.850 ;
        RECT 22.300 38.150 27.700 39.500 ;
        RECT 29.050 38.150 34.450 39.500 ;
        RECT 25.000 35.450 31.750 38.150 ;
        RECT 22.300 34.100 27.700 35.450 ;
        RECT 29.050 34.100 34.450 35.450 ;
        RECT 15.550 32.750 25.000 34.100 ;
        RECT 31.750 32.750 42.550 34.100 ;
        RECT 14.200 31.400 22.300 32.750 ;
        RECT 34.450 31.400 42.550 32.750 ;
        RECT 14.200 30.050 19.600 31.400 ;
        RECT 37.150 30.050 42.550 31.400 ;
        RECT 14.200 28.700 18.250 30.050 ;
        RECT 38.500 28.700 42.550 30.050 ;
        RECT 15.550 27.350 16.900 28.700 ;
        RECT 23.650 27.350 25.000 28.700 ;
        RECT 26.350 27.350 27.700 28.700 ;
        RECT 29.050 27.350 30.400 28.700 ;
        RECT 31.750 27.350 33.100 28.700 ;
        RECT 39.850 27.350 41.200 28.700 ;
        RECT 23.650 24.650 33.100 27.350 ;
        RECT 22.300 23.300 26.350 24.650 ;
        RECT 30.400 23.300 35.800 24.650 ;
        RECT 19.600 21.950 27.700 23.300 ;
        RECT 29.050 21.950 35.800 23.300 ;
        RECT 19.600 20.600 22.300 21.950 ;
        RECT 25.000 20.600 31.750 21.950 ;
        RECT 34.450 20.600 37.150 21.950 ;
        RECT 19.600 19.250 20.950 20.600 ;
        RECT 18.250 17.900 20.950 19.250 ;
        RECT 18.250 16.550 22.300 17.900 ;
        RECT 26.350 16.550 30.400 20.600 ;
        RECT 35.800 19.250 37.150 20.600 ;
        RECT 35.800 17.900 38.500 19.250 ;
        RECT 34.450 16.550 38.500 17.900 ;
        RECT 18.250 11.150 38.500 16.550 ;
        RECT 19.600 8.450 37.150 11.150 ;
        RECT 22.300 7.100 34.450 8.450 ;
        RECT 23.650 5.750 34.450 7.100 ;
  END
END skullfet_inverter
END LIBRARY

